`timescale 1ns / 1ps

`include "neural_network.v"

module neural_network_tb();

    reg [15:0] in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21;
	wire [31:0] out1,out2,out3,out4;

    initial begin 
        $dumpfile("neural_network_tb.vcd");
        $dumpvars(0, neural_network_tb);
    end

    neural_network N1(in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,out1,out2,out3,out4);

    initial begin
        in0 <= 16'b0000_0000_0000_0010;
        in1 <= 16'b0000_0000_0000_0010;
        in2 <= 16'b0000_0000_0000_0010;
        in3 <= 16'b0000_0000_0000_0010;
        in4 <= 16'b0000_0000_0000_0010;
        in5 <= 16'b0000_0000_0000_0010;
        in6 <= 16'b0000_0000_0000_0010;
        in7 <= 16'b0000_0000_0000_0010;
        in8 <= 16'b0000_0000_0000_0010;
        in9 <= 16'b0000_0000_0000_0010;
        in10 <= 16'b0000_0000_0000_0010;
        in11 <= 16'b0000_0000_0000_0010;
        in12 <= 16'b0000_0000_0000_0010;
        in13 <= 16'b0000_0000_0000_0010;
        in14 <= 16'b0000_0000_0000_0010;
        in15 <= 16'b0000_0000_0000_0010;
        in16 <= 16'b0000_0000_0000_0010;
        in17 <= 16'b0000_0000_0000_0010;
        in18 <= 16'b0000_0000_0000_0010;
        in19 <= 16'b0000_0000_0000_0010;
        in20 <= 16'b0000_0000_0000_0010;
        in21 <= 16'b0000_0000_0000_0010;
        
        #1 $display("-----Output1 is %d-----",out1);
        $display("-----Output2 is %d-----",out2);
        $display("-----Output3 is %d-----",out3);
        $display("-----Output4 is %d-----",out4);
        
        #5
        in0 <= 16'b0000_0000_0000_0110;
        in1 <= 16'b0000_0000_0000_1010;
        in2 <= 16'b0000_0000_0000_1010;
        in3 <= 16'b0000_0000_0000_0110;
        in4 <= 16'b0000_0000_0000_0110;
        in5 <= 16'b0000_0000_0000_0110;
        in6 <= 16'b0000_0000_0000_1010;
        in7 <= 16'b0000_0000_0000_1010;
        in8 <= 16'b0000_0000_0000_1110;
        in9 <= 16'b0000_0000_0000_1110;
        in10 <= 16'b0000_0000_0000_1010;
        in11 <= 16'b0000_0000_0000_1010;
        in12 <= 16'b0000_0000_0000_0110;
        in13 <= 16'b0000_0000_0000_0011;
        in14 <= 16'b0000_0000_0000_0011;
        in15 <= 16'b0000_0000_0000_0111;
        in16 <= 16'b0000_0000_0000_0110;
        in17 <= 16'b0000_0000_0000_0010;
        in18 <= 16'b0000_0000_0000_1110;
        in19 <= 16'b0000_0000_0000_1010;
        in20 <= 16'b0000_0000_0000_1010;
        in21 <= 16'b0000_0000_0000_0110;
        
        #1 $display("\n-----Output1 is %d-----",out1);
        $display("-----Output2 is %d-----",out2);
        $display("-----Output3 is %d-----",out3);
        $display("-----Output4 is %d-----",out4);
        
        #5
        in0 <= 16'b0000_0000_0001_0110;
        in1 <= 16'b0000_0000_0000_1010;
        in2 <= 16'b0000_0000_0000_1010;
        in3 <= 16'b0000_0000_0000_0110;
        in4 <= 16'b0000_0000_0000_0110;
        in5 <= 16'b0000_0000_0000_0110;
        in6 <= 16'b0000_0000_0000_1010;
        in7 <= 16'b0000_0000_0000_1010;
        in8 <= 16'b0000_0000_0000_1110;
        in9 <= 16'b0000_0000_0000_1110;
        in10 <= 16'b0000_0000_0000_1010;
        in11 <= 16'b0000_0000_0000_1010;
        in12 <= 16'b0000_0000_0000_0110;
        in13 <= 16'b0000_0000_0000_0011;
        in14 <= 16'b0000_0000_0000_0011;
        in15 <= 16'b0000_0000_0000_0111;
        in16 <= 16'b0000_0000_0000_0110;
        in17 <= 16'b0000_0000_0000_0010;
        in18 <= 16'b0000_0000_0000_1110;
        in19 <= 16'b0000_0000_0000_1010;
        in20 <= 16'b0000_0000_0000_1010;
        in21 <= 16'b0000_0000_0000_0110;
        
        #1 $display("\n-----Output1 is %d-----",out1);
        $display("-----Output2 is %d-----",out2);
        $display("-----Output3 is %d-----",out3);
        $display("-----Output4 is %d-----",out4);
        
        #1 $finish;
    end
endmodule